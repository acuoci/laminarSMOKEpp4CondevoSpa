! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: POLIMI_TOT_NOx_1407.CKT
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 1/20/2017

THERMO ALL
270.   1000.   3500. 
CH4                     C   1H   4          G    300.00   3500.00 1070.00      1
-2.82321418e-01 1.42739336e-02-6.77628877e-06 1.55380951e-09-1.39473841e-13    2
-9.36383584e+03 2.03507025e+01 2.85765313e+00 2.53571099e-03 9.67916347e-06    3
-8.69880871e-09 2.25599771e-12-1.00357904e+04 4.98969391e+00                   4
O2                      O   2               G    300.00   3500.00  760.00      1
 2.81750647e+00 2.49838008e-03-1.52493522e-06 4.50547610e-10-4.87702795e-14    2
-9.31713391e+02 7.94729338e+00 3.46035081e+00-8.85011180e-04 5.15281069e-06    3
-5.40712424e-09 1.87809546e-12-1.02942573e+03 5.02236122e+00                   4
CO2                     C   1O   2          G    300.00   3500.00 1620.00      1
 5.07830985e+00 2.05366041e-03-5.94311264e-07 5.38675127e-11 1.66346859e-15    2
-4.92442103e+04-4.47815291e+00 2.44892797e+00 8.54596135e-03-6.60570102e-06    3
 2.52769046e-09-3.80099332e-13-4.83922906e+04 9.47557732e+00                   4
CO                      C   1O   1          G    300.00   3500.00 1000.00      1
 2.68595014e+00 2.12486373e-03-1.04548609e-06 2.45538865e-10-2.22550982e-14    2
-1.41423615e+04 7.96579427e+00 3.81890943e+00-2.40697344e-03 5.75226967e-06    3
-4.28629830e-09 1.11070419e-12-1.43689533e+04 2.49992059e+00                   4
H2O                     H   2O   1          G    300.00   3500.00 1590.00      1
 2.30940463e+00 3.65433887e-03-1.22983871e-06 2.11931684e-10-1.50333493e-14    2
-2.97294901e+04 8.92765177e+00 4.03530937e+00-6.87559834e-04 2.86629215e-06    3
-1.50552360e-09 2.55006790e-13-3.02783278e+04-1.99201641e-01                   4
H2                      H   2               G    300.00   3500.00  750.00      1
 3.73110903e+00-8.86706228e-04 1.12286898e-06-3.74349786e-10 4.17963679e-14    2
-1.08851547e+03-5.35285858e+00 3.08866001e+00 2.53968852e-03-5.72992051e-06    3
 5.71701866e-09-1.98865978e-12-9.92148122e+02-2.43823451e+00                   4
H                       H   1               G    300.00   3500.00 1800.00      1
 2.50000000e+00-3.95459854e-15 2.96893838e-18-9.33318862e-22 1.04354326e-25    2
 2.54716200e+04-4.60117600e-01 2.50000000e+00 1.70660813e-16-4.68777753e-19    3
 3.39909334e-22-7.24829229e-26 2.54716200e+04-4.60117600e-01                   4
O                       O   1               G    300.00   3500.00  950.00      1
 2.57318360e+00-8.95609973e-05 4.05096293e-08-8.39812642e-12 9.43621954e-16    2
 2.92191409e+04 4.74952023e+00 2.95200330e+00-1.68459131e-03 2.55897855e-06    3
-1.77574473e-09 4.66034835e-13 2.91471652e+04 2.94136507e+00                   4
OH                      H   1O   1          G    300.00   3500.00  880.00      1
 3.62538437e+00-5.02165284e-04 8.36958465e-07-2.95714532e-10 3.30350487e-14    2
 3.41380110e+03 1.55419439e+00 3.37995108e+00 6.13440537e-04-1.06464237e-06    3
 1.14489216e-09-3.76228216e-13 3.45699735e+03 2.70689353e+00                   4
HO2                     H   1O   2          G    300.00   3500.00 1540.00      1
 4.16318067e+00 1.99798265e-03-4.89192085e-07 7.71153169e-11-7.30772101e-15    2
 4.41348946e+01 2.95517985e+00 2.85241381e+00 5.40257188e-03-3.80535043e-06    3
 1.51268170e-09-2.40354212e-13 4.47851086e+02 9.84483831e+00                   4
CH2                     C   1H   2          G    300.00   3500.00  900.00      1
 3.24505871e+00 2.75395076e-03-7.68471345e-07 8.23040044e-11-1.89900259e-15    2
 4.54794580e+04 4.28187007e+00 3.99717917e+00-5.88806836e-04 4.80279131e-06    3
-4.04455722e-09 1.14445134e-12 4.53440763e+04 7.32567425e-01                   4
CH2S                    C   1H   2          G    300.00   3500.00  900.00      1
 2.57518274e+00 4.11179660e-03-1.68232436e-06 3.44404950e-10-2.93085970e-14    2
 5.01958500e+04 6.99914505e+00 4.62572655e+00-5.00173142e-03 1.35068890e-05    3
-1.09068642e-08 3.09604395e-12 4.98267521e+04-2.67749713e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1270.00      1
 2.57723974e+00 6.62601164e-03-2.54906392e-06 4.67320141e-10-3.34867663e-14    2
 1.65488693e+04 6.94195966e+00 3.53327401e+00 3.61488008e-03 1.00739068e-06    3
-1.39958516e-09 3.34014278e-13 1.63060366e+04 2.10113860e+00                   4
HCO                     C   1H   1O   1     G    300.00   3500.00  920.00      1
 2.44772077e+00 5.65570556e-03-3.01329556e-06 7.57702525e-10-7.26129632e-14    2
 4.31149160e+03 1.15871953e+01 3.74218864e+00 2.75843940e-05 6.16298894e-06    3
-5.89177900e-09 1.73431136e-12 4.07330951e+03 5.45007089e+00                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  930.00      1
 1.06639253e+00 1.06960337e-02-5.54447373e-06 1.36053696e-09-1.28442555e-13    2
-1.46324373e+04 1.74071779e+01 3.13463322e+00 1.80037481e-03 8.80336319e-06    3
-8.92465079e-09 2.63639286e-12-1.50171301e+04 7.57920579e+00                   4
CH3OO                   C   1H   3O   2     G    300.00   3500.00 1300.00      1
 3.46521970e+00 1.23938518e-02-5.59614682e-06 1.22616716e-09-1.06238815e-13    2
 6.86982281e+02 1.04298931e+01 4.30117244e+00 9.82168948e-03-2.62826727e-06    3
-2.95822350e-10 1.86451475e-13 4.69634569e+02 6.17758023e+00                   4
C2H4                    C   2H   4          G    300.00   3500.00 1800.00      1
 4.49333672e+00 1.00335105e-02-3.62601388e-06 5.97613541e-10-3.65481279e-14    2
 3.93220822e+03-3.35192021e+00 2.66161697e-01 1.94272328e-02-1.14541158e-05    3
 3.49691054e-09-4.39228267e-13 5.45399123e+03 1.95264329e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00  700.00      1
-1.10489358e+00 2.43511913e-02-1.39613152e-05 3.89870297e-09-4.17285120e-13    2
 1.35030749e+04 3.00146907e+01 4.99501829e+00-1.05054480e-02 6.07314832e-05    3
-6.72372955e-08 2.49884286e-11 1.26490872e+04 2.76182769e+00                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1800.00      1
 7.44900313e+00 1.01177830e-03 3.02918166e-07-2.13909391e-10 2.81815209e-14    2
 1.86458955e+04-1.30987733e+01 4.44514163e+00 7.68702607e-03-5.25978830e-06    3
 1.84635226e-09-2.57965931e-13 1.97272856e+04 3.15875175e+00                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1410.00      1
 6.03578795e+00 5.81722421e-03-1.93206512e-06 2.83140053e-10-1.50051611e-14    2
-8.58422380e+03-7.64505060e+00 2.49197065e+00 1.58706066e-02-1.26271528e-05    3
 5.33991909e-09-9.11597189e-13-7.58486732e+03 1.06694385e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1030.00      1
 3.66502520e+00 1.44768244e-02-7.23266377e-06 1.70580456e-09-1.56345856e-13    2
-3.68579206e+01 5.92341848e+00 2.15742064e-01 2.78720987e-02-2.67403448e-05    3
 1.43321353e-08-3.22098925e-12 6.73694407e+02 2.26661724e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00  700.00      1
 7.05094232e-01 1.53761148e-02-8.91788177e-06 2.51340904e-09-2.70561650e-13    2
 3.36189510e+04 1.96531878e+01 2.74606707e+00 3.71341285e-03 1.60736223e-05    3
-2.12880234e-08 8.22994995e-12 3.33332148e+04 1.05346375e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  970.00      1
 4.61193612e+00 5.01498203e-03-1.65253693e-06 2.49922529e-10-1.30568633e-14    2
 2.56043843e+04-3.75517098e+00 1.83812159e+00 1.64533925e-02-1.93408005e-05    3
 1.24068047e-08-3.14627392e-12 2.61425043e+04 9.54239254e+00                   4
N2                      N   2               G    300.00   3500.00 1050.00      1
 2.71287897e+00 1.90359754e-03-8.54297558e-07 1.84170938e-10-1.54715989e-14    2
-8.40225273e+02 7.15926558e+00 3.85321337e+00-2.44053350e-03 5.35160392e-06    3
-3.75608397e-09 9.22684332e-13-1.07969550e+03 1.60217419e+00                   4
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
!NOx MODULE (from Burcat http://garfield.chem.elte.hu/Burcat/THERM.DAT)
!+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NO                RUS 89N   1O   1    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.26071234E+00 1.19101135E-03-4.29122646E-07 6.94481463E-11-4.03295681E-15    2
 9.92143132E+03 6.36900518E+00 4.21859896E+00-4.63988124E-03 1.10443049E-05    3
-9.34055507E-09 2.80554874E-12 9.84509964E+03 2.28061001E+00 1.09770882E+04    4
N2O               L 7/88N   2O   1    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 0.48230729E+01 0.26270251E-02-0.95850872E-06 0.16000712E-09-0.97752302E-14    2
 0.80734047E+04-0.22017208E+01 0.22571502E+01 0.11304728E-01-0.13671319E-04    3
 0.96819803E-08-0.29307182E-11 0.87417746E+04 0.10757992E+02 0.98141682E+04    4
NO2               L 7/88N   1O   2    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 0.48847540E+01 0.21723955E-02-0.82806909E-06 0.15747510E-09-0.10510895E-13    2
 0.23164982E+04-0.11741695E+00 0.39440312E+01-0.15854290E-02 0.16657812E-04    3
-0.20475426E-07 0.78350564E-11 0.28966180E+04 0.63119919E+01 0.41124701E+04    4
HNO               ATcT/AH  1.N  1.O  1.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.16598124E+00 2.99958892E-03-3.94376786E-07-3.85344089E-11 7.07602668E-15    2
 1.17726311E+04 7.64511172E+00 4.53525574E+00-5.68543377E-03 1.85198540E-05    3
-1.71881225E-08 5.55818157E-12 1.16183003E+04 1.74315886E+00 1.28500657E+04    4
HNO2              ATcT3EH   1N   1O   2    0G    200.00   6000.00 1000.00      1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 4.66358504E+00 4.89854351E-03-1.79694193E-06 2.94420361E-10-1.78235577E-14    2
-7.25216334E+03-3.06053640E-02 4.03779347E+00-4.46123109E-03 3.19440815E-05    3
-3.79359490E-08 1.44570885E-11-6.53088236E+03 5.90620097E+00-5.31122753E+03    4
HONO              ATcT3EH   1N   1O   2    0G    200.00   6000.00 1000.00      1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 5.79144641E+00 3.64630732E-03-1.29112765E-06 2.06498233E-10-1.22138679E-14    2
-1.15974343E+04-4.07145349E+00 3.16416438E+00 8.50517773E-03 5.48561573E-07    3
-8.27656474E-09 4.39957151E-12-1.07744086E+04 1.00231941E+01-9.46242812E+03    4
HONO2             T 8/03H  1.N  1.O  3.   0.G   200.000  6000.000 1000.        1 ! HNO3 in Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 8.03098942E+00 4.46958589E-03-1.72459491E-06 2.91556153E-10-1.80102702E-14    2
-1.93138183E+04-1.62616537E+01 1.69329154E+00 1.90167702E-02-8.25176697E-06    3
-6.06113827E-09 4.65236978E-12-1.74198909E+04 1.71839838E+01-1.61524852E+04    4
N2H2      2/13/19       N   2H   2          G   300.000  5000.000 1380.000     1 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 4.14686796E+00 4.81612315E-03-1.62748817E-06 2.50556098E-10-1.44494188E-14    2
 2.33444055E+04 5.34122740E-01 2.55589425E+00 6.54339081E-03-8.81947855E-07    3
-1.15971304E-09 3.97442230E-13 2.41085081E+04 9.80504705E+00                   4
H2NN Isodiazene   T 9/11N  2.H  2.   0.   0.G   200.000  6000.000 1000.        1 ! Is 'N2H2 Isodiazene' in Burcat database
 3.05903670E+00 6.18382347E-03-2.22171165E-06 3.58539206E-10-2.14532905E-14    2
 3.48530149E+04 6.69893515E+00 4.53204001E+00-7.32418578E-03 3.00803713E-05    3
-3.04000551E-08 1.04700639E-11 3.49580003E+04 1.51074195E+00 3.61943157E+04    4
HNNO      5/30/18 THERM N  2.H  1.O  1    0.G   300.000  5000.000 1790.000    61 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 2.15594002E+06-4.13111192E+03 2.65627771E+00-6.70395293E-04 5.57827338E-08    2
-8.03468100E+08-1.18702032E+07-8.96779017E-01 3.69714359E-02-4.80099825E-05    3
 2.62274393E-08-5.11382966E-12 2.68675048E+04 2.64521806E+01                   4
NH2NO     5/30/18 THERM N  2.H  2.O  1    0.G   300.000  5000.000 1371.000    61 ! Dean AM Bozzelli JW (Gardiner WC) Gas Phase Combustion Chemistry, Springer 2000.
 7.93898100E+00 5.21842622E-03-2.12493130E-06 3.53331059E-10-2.12447889E-14    2
 5.42322972E+03-1.84299492E+01 1.85914077E+00 1.68525394E-02-9.37240888E-06    3
 1.71380329E-09 4.84625807E-14 7.78108234E+03 1.51172833E+01                   4
HNOH trans & Equ  T11/11H  2.N  1.O  1.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.98321933E+00 4.88846374E-03-1.65086637E-06 2.55371446E-10-1.48308561E-14    2
 1.05780106E+04 3.62582838E+00 3.95608248E+00-3.02611020E-03 2.56874396E-05    3
-3.15645120E-08 1.24084574E-11 1.09199790E+04 5.55950983E+00 1.21354115E+04    4
NH2OH             ATcT/AN  1.H  3.O  1.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.88112502E+00 8.15708448E-03-2.82615576E-06 4.37930933E-10-2.52724604E-14    2
-6.86018419E+03 3.79156136E+00 3.21016092E+00 6.19671676E-03 1.10594948E-05    3
-1.96668262E-08 8.82516590E-12-6.58148481E+03 7.93293571E+00-5.28593988E+03    4
NH3               ATcT3EH   3N   1    0    0G    200.00   4000.00 1000.00      1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 2.36074311E+00 6.31850146E-03-2.28966806E-06 4.11767411E-10-2.90836787E-14    2
-6.41596473E+03 8.02154329E+00 4.14027871E+00-3.58489142E-03 1.89475904E-05    3
-1.98833970E-08 7.15267961E-12-6.68545158E+03-1.66754883E-02-5.47888720E+03    4
N2H4 HYDRAZINE    L 5/90N   2H   4    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 4.93957357E+00 8.75017187E-03-2.99399058E-06 4.67278418E-10-2.73068599E-14    2
 9.28265548E+03-2.69439772E+00 3.83472149E+00-6.49129555E-04 3.76848463E-05    3
-5.00709182E-08 2.03362064E-11 1.00893925E+04 5.75272030E+00 1.14474575E+04    4
N                 L 6/88N   1    0    0    0G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 0.24159429E+01 0.17489065E-03-0.11902369E-06 0.30226244E-10-0.20360983E-14    2
 0.56133775E+05 0.46496095E+01 0.25000000E+01 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.56104638E+05 0.41939088E+01 0.56850013E+05    4
NO3               ATcT/AN  1.O  3.   0.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 7.48347702E+00 2.57772064E-03-1.00945831E-06 1.72314063E-10-1.07154008E-14    2
 6.12990474E+03-1.41618136E+01 2.17359330E+00 1.04902685E-02 1.10472669E-05    3
-2.81561867E-08 1.36583960E-11 7.81290905E+03 1.46022090E+01 8.97563416E+03    4
NH                ATcT/AN  1.H  1.   0.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 2.78372644E+00 1.32985888E-03-4.24785573E-07 7.83494442E-11-5.50451310E-15    2
 4.23461945E+04 5.74084863E+00 3.49295037E+00 3.11795720E-04-1.48906628E-06    3
 2.48167402E-09-1.03570916E-12 4.21059722E+04 1.84834973E+00 4.31525130E+04    4
NNH               T 8/11N  2.H  1.   0.   0.G   200.000  6000.000 1000.        1 ! N2H in Burcat database http://garfield.chem.elte.hu/Burcat/THERM.DAT
 3.42744423E+00 3.23295234E-03-1.17296299E-06 1.90508356E-10-1.14491506E-14    2
 2.87676026E+04 6.39209233E+00 4.25474632E+00-3.45098298E-03 1.37788699E-05    3
-1.33263744E-08 4.41023397E-12 2.87932080E+04 3.28551762E+00 3.00058572E+04    4
NH2  AMIDOGEN RAD IU3/03N  1.H  2.   0.   0.G   200.000  3000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 2.59263049E+00 3.47683597E-03-1.08271624E-06 1.49342558E-10-5.75241187E-15    2
 2.15737320E+04 7.90565351E+00 4.19198016E+00-2.04602827E-03 6.67756134E-06    3
-5.24907235E-09 1.55589948E-12 2.11863286E+04-9.04785244E-02 2.23945849E+04    4
H2NO  RADICAL     T09/09N  1.H  2.O  1.   0.G   200.000  6000.000 1000.        1 ! Glarborg, P. et al. Progr Energy Combust Sci, 67, 31-68. (2018)
 3.75555914E+00 5.16219354E-03-1.76387387E-06 2.75052692E-10-1.60643143E-14    2
 6.51826177E+03 4.30933053E+00 3.93201139E+00-1.64028165E-04 1.39161409E-05    3
-1.62747853E-08 6.00352834E-12 6.71178975E+03 4.58837038E+00 7.97044877E+03    4
N2H3   Rad.       T 7/11N  2.H  3.   0.   0.G   200.000  6000.000 1000.        1 ! E. Goos, A. Burcat and B. Ruscic http://garfield.chem.elte.hu/Burcat/THERM.DAT
 4.04483566E+00 7.31130186E-03-2.47625799E-06 3.83733021E-10-2.23107573E-14    2
 2.53241420E+04 2.88423392E+00 3.42125505E+00 1.34901590E-03 2.23459071E-05    3
-2.99727732E-08 1.20978970E-11 2.58198956E+04 7.83176309E+00 2.70438066E+04    4
END
